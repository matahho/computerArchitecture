module adder(a, b,o);
    input [31:0] a, b;
    output [31:0]o;

    
    assign o = a + b;
endmodule
